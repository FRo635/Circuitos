module demux(d0, s0, s1, y0, y1, y2, y3)

    input = d0, s0, s1
    output = y0, y1, y2, y3