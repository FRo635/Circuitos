module mux(s0, s1, s2, s3, y)

    input = s0, s1, s2, s3

    output reg Y;

    assign Y  =


endmodule