module demux(s0, s1, y0, y1, y2, y3)